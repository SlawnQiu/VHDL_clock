LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY BEEPCTRL IS
PORT(
	CLK : IN STD_LOGIC;
	SW1, START1, START2 : IN STD_LOGIC;
	BEEPER : OUT STD_LOGIC
	);
END ENTITY;

ARCHITECTURE BEHAV OF BEEPCTRL IS

TYPE MODE IS (UP, DOWN);
SIGNAL STATE : MODE := DOWN;
SIGNAL TMP, TMP1, TMP2, SW1_DROP, START1_RISE, START2_RISE : STD_LOGIC;
BEGIN

PROCESS(CLK)
BEGIN
IF CLK'EVENT AND CLK='1' THEN
	TMP <= SW1;
END IF;
END PROCESS;
SW1_DROP <= '0' WHEN (SW1='0' AND TMP ='1') ELSE '1';

PROCESS(CLK)
BEGIN
IF CLK'EVENT AND CLK='1' THEN
	TMP1 <= START1;
END IF;
END PROCESS;
START1_RISE <= '1' WHEN (START1='1' AND TMP1 ='0') ELSE '0';

PROCESS(CLK)
BEGIN
IF CLK'EVENT AND CLK='1' THEN
	TMP2 <= START2;
END IF;
END PROCESS;
START2_RISE <= '1' WHEN (START2='1' AND TMP2 ='0') ELSE '0';

PROCESS(CLK, SW1_DROP, START1_RISE, START2_RISE)
BEGIN
	IF RISING_EDGE(CLK) THEN
		CASE STATE IS
			WHEN UP =>
				IF SW1_DROP = '0' THEN
					STATE <= DOWN;
				END IF;
			WHEN DOWN =>
				IF START1_RISE = '1' OR START2_RISE = '1' THEN
					STATE <= UP;
				END IF;
		END CASE;
	END IF;
END PROCESS;

PROCESS(CLK)		--OUTPUT
BEGIN
IF RISING_EDGE(CLK) THEN
	CASE STATE IS
		WHEN UP =>
			BEEPER <= '1';
		WHEN DOWN =>
			BEEPER <= '0';
		WHEN OTHERS => NULL;
	END CASE;
END IF;
END PROCESS;

END BEHAV;