LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
ENTITY CLK_GEN IS
	PORT(
		CLKIN: IN STD_LOGIC;
		OCLK1K, OCLK2HZ, OCLK1HZ: OUT STD_LOGIC
		);
END CLK_GEN;

ARCHITECTURE FLOW OF CLK_GEN IS
SIGNAL	CLK1M: STD_LOGIC;
SIGNAL	TIME50: INTEGER RANGE 0 TO 49;
SIGNAL	CLK1K: STD_LOGIC;
SIGNAL	TIME1K: INTEGER RANGE 0 TO 999;
SIGNAL	CLK2HZ: STD_LOGIC;
SIGNAL	TIME500: INTEGER RANGE 0 TO 499;
SIGNAL	CLK1HZ: STD_LOGIC;
SIGNAL	TIME2: INTEGER RANGE 0 TO 1;


BEGIN


PROCESS(CLKIN) --1/50
BEGIN
IF CLKIN 'EVENT AND CLKIN = '1' THEN
	TIME50 <= TIME50 + 1;
	IF TIME50 = 49 THEN
		CLK1M <= '1';
		TIME50 <= 0;
	ELSE
		CLK1M <= '0';
	END IF;
END IF;
END PROCESS;

PROCESS(CLK1M) --1/50000
BEGIN
IF CLK1M 'EVENT AND CLK1M = '1' THEN
	TIME1K <= TIME1K + 1;
	IF TIME1K = 999 THEN
		CLK1K <= '1';
		TIME1K <= 0;
	ELSE
		CLK1K <= '0';
	END IF;
END IF;
END PROCESS;

PROCESS(CLK1K)
BEGIN
OCLK1K <= CLK1K;
END PROCESS;

PROCESS(CLK1K) --1/25000000
BEGIN
IF CLK1K 'EVENT AND CLK1K = '1' THEN
	TIME500 <= TIME500 + 1;
	IF TIME500 = 499 THEN
		CLK2HZ <= '1';
		TIME500 <= 0;
	ELSE
		CLK2HZ <= '0';
	END IF;
END IF;
END PROCESS;

PROCESS(CLK2HZ)
BEGIN
OCLK2HZ <= CLK2HZ;
END PROCESS;

PROCESS(CLK2HZ) --1/25000000
BEGIN
IF CLK2HZ 'EVENT AND CLK2HZ = '1' THEN
	TIME2 <= TIME2 + 1;
	IF TIME2 = 1 THEN
		CLK1HZ <= '1';
		TIME2 <= 0;
	ELSE
		CLK1HZ <= '0';
	END IF;
END IF;
END PROCESS;

PROCESS(CLK1HZ)
BEGIN
OCLK1HZ <= CLK1HZ;
END PROCESS;

END FLOW;