LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
ENTITY COMPARATOR IS
	PORT(
			CLK, EN : IN STD_LOGIC;
			BEEP : OUT STD_LOGIC;
			I2SEC0, I2SEC1, I2MIN0, I2MIN1, I2HR0, I2HR1 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			I1SEC0, I1SEC1, I1MIN0, I1MIN1, I1HR0, I1HR1 : IN STD_LOGIC_VECTOR(3 DOWNTO 0)
		);
END ENTITY;

ARCHITECTURE BEHAV OF COMPARATOR IS
BEGIN
PROCESS(CLK)
BEGIN
IF RISING_EDGE(CLK) THEN
	IF EN = '1' THEN
		IF I1HR0 = I2HR0 AND I1HR1 = I2HR1 AND I1SEC0 = I2SEC0 AND I1SEC1 = I2SEC1 AND I1MIN0 = I2MIN0 AND I1MIN1 = I2MIN1 THEN
			BEEP <= '1';
		ELSE
			BEEP <= '0';
		END IF;
	ELSE
		BEEP <= '0';
	END IF;
END IF;
END PROCESS;

END BEHAV;