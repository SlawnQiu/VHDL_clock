LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
ENTITY CLK_GEN IS
	PORT(
		CLKIN: IN STD_LOGIC;
		OCLK1K, OCLK2HZ, OCLK1HZ: OUT STD_LOGIC
		);
END CLK_GEN;

ARCHITECTURE FLOW OF CLK_GEN IS
SIGNAL COUNT5W: INTEGER RANGE 1 TO 50000;
SIGNAL COUNT25M: INTEGER RANGE 1 TO 25000000;
SIGNAL COUNT50M: INTEGER RANGE 1 TO 50000000;

BEGIN

PROCESS(CLKIN)			--GENERATE 1KHZ
BEGIN
	IF RISING_EDGE(CLKIN) THEN
		COUNT5W <= COUNT5W + 1;
		IF(COUNT5W >= 25000)THEN
			OCLK1K <= '1';
		ELSE
			OCLK1K <= '0';
		END IF;
		IF COUNT5W = 50000 THEN
			COUNT5W <= 1;
		END IF;
	END IF;
END PROCESS;

PROCESS(CLKIN)			--GENERATE 2HZ
BEGIN
	IF RISING_EDGE(CLKIN) THEN
		COUNT25M <= COUNT25M + 1;
		IF(COUNT25M >= 12500000)THEN
			OCLK2HZ <= '1';
		ELSE
			OCLK2HZ <= '0';
		END IF;
		IF COUNT25M = 25000000 THEN
			COUNT25M <= 1;
		END IF;
	END IF;
END PROCESS;


PROCESS(CLKIN)			--GENERATE 1HZ
BEGIN
	IF RISING_EDGE(CLKIN) THEN
		COUNT50M <= COUNT50M + 1;
		IF(COUNT50M >= 25000000)THEN
			OCLK1HZ <= '1';
		ELSE
			OCLK1HZ <= '0';
		END IF;
		IF COUNT50M = 50000000 THEN
			COUNT50M <= 1;
		END IF;
	END IF;
END PROCESS;

END FLOW;